/*
=============================================================
    Owners      : Everyone (Grecia, Manuel, Emmanuel, German)
    Last update    : 03 Jul 2023 by German
=============================================================            
*/

package ram_env_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

    `include "port1_agent/ram_port1_sequence_item.svh"
    // `include "port1_agent/ram_port1_monitor.svh"
    // `include "port1_agent/ram_port1_scb.svh"
    // `include "port1_agent/ram_port1_subs.svh"
    `include "port1_agent/ram_port1_sequencer.svh"
    `include "port1_agent/ram_port1_driver.svh"
    `include "port1_agent/ram_port1_agent.svh"
    
	// `include "ram_env.svh"

endpackage