`define ADDR_WIDTH 'd8
`define DATA_WIDTH 'd32 
`define clk0_period 10
`define clk1_period 10